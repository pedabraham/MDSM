library IEEE;
